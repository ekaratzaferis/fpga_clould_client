`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   17:35:35 10/23/2014
// Design Name:   dvi_drawer
// Module Name:   C:/VHDL/fpga_client_v2/tb_dvi_drawer.v
// Project Name:  fpga_client_v2
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: dvi_drawer
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module tb_dvi_drawer;

	// Inputs
	reg pixel_clock;
	reg new_frame;
	reg new_line;
	reg ram_ack;
	reg ram_init;
	reg [6143:0] read_data;

	// Outputs
	wire ask_data;
	wire [7:0] R;
	wire [7:0] G;
	wire [7:0] B;

	// Instantiate the Unit Under Test (UUT)
	dvi_drawer uut (
		.pixel_clock(pixel_clock), 
		.new_frame(new_frame), 
		.new_line(new_line), 
		.ask_data(ask_data), 
		.ram_init(ram_init), 
		.R(R), 
		.G(G), 
		.B(B), 
		.ram_ack(ram_ack), 
		.read_data(read_data)
	);

	initial begin
		// Initialize Inputs
		pixel_clock = 0;
		new_frame = 0;
		new_line = 0;
		ram_init = 0;
		ram_ack = 0;
		read_data = 0;

		// Wait 100 ns for global reset to finish
		#100;
		read_data <= 6144'h012345678955667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677889900112233445566778899001122334455667788990011223344556677;

		@(posedge pixel_clock);
		new_frame = 1;
		new_line = 1;
		ram_init = 1;
		@(posedge pixel_clock);
		new_frame = 0;
		new_line = 0;
		
		#240;
		@(posedge pixel_clock);
		ram_ack = 1;
		@(posedge pixel_clock);
		ram_ack = 0;
		
		#20600;
		@(posedge pixel_clock);
		new_line = 1;
		@(posedge pixel_clock);
		new_line = 0;
		
		#10000000;
		@(posedge pixel_clock);
		new_frame = 1;
		@(posedge pixel_clock);
		new_frame = 0;
		
	end
      
	always begin	
		#10;
		pixel_clock = ~pixel_clock;
	end
      
endmodule

